module exception_pchandling(output  logic [31:0] MoveR14PC_D);

	assign MoveR14PC_D = 32'b1110_000_1101_0_0000_1110_00000000_1111;

endmodule 