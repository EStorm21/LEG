/*
   LEG Processor for Education
   Copyright (C) 2016  Max Waugaman

   This program is free software: you can redistribute it and/or modify
   it under the terms of the GNU General Public License as published by
   the Free Software Foundation, either version 3 of the License, or
   (at your option) any later version.

   This program is distributed in the hope that it will be useful,
   but WITHOUT ANY WARRANTY; without even the implied warranty of
   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
   GNU General Public License for more details.

   You should have received a copy of the GNU General Public License
   along with this program.  If not, see <http://www.gnu.org/licenses/>.
*/

module tlb #(parameter tbits = 16, parameter size = 16, 
parameter tlb_word_size = tbits   + 1        + 1          + 2  + 4      + 1)
//                        phystag + cachable + bufferable + AP + Domain + valid
(
    input logic clk, reset, enable, we, // Clock
    input logic [tbits-1:0] VirtTag,
    inout logic [tlb_word_size-1:0] TableEntry, // Physical Tag to write data into TLB
    output logic PAReady
);

/***** Brief Description *******
 * First Created by Max Waugaman 2015
 *
 * tlb uses a CAM connected to a match RAM to perform virtual to physical
 * address translation. The current addressing policy uses an index of the
 * virtual address to determine the location of the entry in the CAM and RAM.
 ******************************/


// RAM signals
tri [tlb_word_size-1:0] RData;
logic                     RRead ;

// CAM signals
logic [$size(VirtTag) - 1:0] CData ;
logic [  $clog2(size) - 1:0] CAdr  ;
logic                        CRead ;

// Shared Signals
logic [size - 1:0] Match;
logic [size - 1:0] WriteMatch; // TODO: Remove, make match < 1 cycle
logic [size - 1:0] CamMatch; // TODO: Remove, make match < 1 cycle

// Valid signal for controller
logic valid;

// The match signal is not generated by the CAM in time for a write to the RAM
// In a physical implementation, for subcycle TLB acesses, the CAM would have 
// to generate the Match signal in less than one cycle. Here, we create a 
// separate write address to avoid this problem and use simple memory in 
// the match_ram and tlb_controller.
onehot16 onehotMatch(CAdr, WriteMatch);
mux2 #(size) matchMux(CamMatch, WriteMatch, we, Match);

cam #(tbits, size) 
tlb_cam(clk, reset, enable, CRead, we, CAdr, CData, CamMatch);

match_ram #(tlb_word_size, size) 
tlb_ram(clk, reset, enable, RRead, we, Match, RData);

tlb_controller #(size, tbits) tc(.*);

assign valid = TableEntry[0];
assign RData = we ? TableEntry : 'bz;
assign CData = VirtTag;
assign TableEntry = !we ? RData : 'bz;
assign Miss = ~(|Match) | ~valid;

endmodule
