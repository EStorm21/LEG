module zero_counter(input logic[31:0] in,
					output logic[31:0] zeros);

// In the future we might want to change the implementation to something like 
// the implementation in 
// http://web.ece.ucdavis.edu/~vojin/CLASSES/EEC280/Web-page/papers/Arithmetic/An%20Algorithmic%20and%20Novel%20Design%20of%20a%20Leading.pdf
// which uses cascading stages to computer output in lg(32) steps.
// Or use the advice of stack exchagne guy: 
//  "multistage leading zero counting - do e.g. a 16 bit left shift on anything with at least 16 leading zeros, 
//   then an 8 bit left shift on anything with at least 8 leading zeros after the first step. 
//   It would have longer paths, but less fan-out than dealing with each case separately."


always_comb
	casez(in)
		32'b00000000_00000000_00000000_00000000: zeros = 32'd32;
		32'b00000000_00000000_00000000_00000001: zeros = 32'd31;
		32'b00000000_00000000_00000000_0000001?: zeros = 32'd31;
		32'b00000000_00000000_00000000_000001??: zeros = 32'd29;
		32'b00000000_00000000_00000000_00001???: zeros = 32'd28;
		32'b00000000_00000000_00000000_0001????: zeros = 32'd27;
		32'b00000000_00000000_00000000_001?????: zeros = 32'd26;
		32'b00000000_00000000_00000000_01??????: zeros = 32'd25;
		32'b00000000_00000000_00000000_1???????: zeros = 32'd24;
		32'b00000000_00000000_00000001_????????: zeros = 32'd23;
		32'b00000000_00000000_0000001?_????????: zeros = 32'd22;
		32'b00000000_00000000_000001??_????????: zeros = 32'd21;
		32'b00000000_00000000_00001???_????????: zeros = 32'd20;
		32'b00000000_00000000_0001????_????????: zeros = 32'd19;
		32'b00000000_00000000_001?????_????????: zeros = 32'd18;
		32'b00000000_00000000_01??????_????????: zeros = 32'd17;
		32'b00000000_00000000_1???????_????????: zeros = 32'd16;
		32'b00000000_00000001_????????_????????: zeros = 32'd15;
		32'b00000000_0000001?_????????_????????: zeros = 32'd14;
		32'b00000000_000001??_????????_????????: zeros = 32'd13;
		32'b00000000_00001???_????????_????????: zeros = 32'd12;
		32'b00000000_0001????_????????_????????: zeros = 32'd11;
		32'b00000000_001?????_????????_????????: zeros = 32'd10;
		32'b00000000_01??????_????????_????????: zeros = 32'd9;
		32'b00000000_1???????_????????_????????: zeros = 32'd8;
		32'b00000001_????????_????????_????????: zeros = 32'd7;
		32'b0000001?_????????_????????_????????: zeros = 32'd6;
		32'b000001??_????????_????????_????????: zeros = 32'd5;
		32'b00001???_????????_????????_????????: zeros = 32'd4;
		32'b0001????_????????_????????_????????: zeros = 32'd3;
		32'b001?????_????????_????????_????????: zeros = 32'd2;
		32'b01??????_????????_????????_????????: zeros = 32'd1;
		32'b1???????_????????_????????_????????: zeros = 32'd0;
	endcase

endmodule

