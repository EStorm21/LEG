/*
   LEG Processor for Education
   Copyright (C) 2016  Max Waugaman

   This program is free software: you can redistribute it and/or modify
   it under the terms of the GNU General Public License as published by
   the Free Software Foundation, either version 3 of the License, or
   (at your option) any later version.

   This program is distributed in the hope that it will be useful,
   but WITHOUT ANY WARRANTY; without even the implied warranty of
   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
   GNU General Public License for more details.

   You should have received a copy of the GNU General Public License
   along with this program.  If not, see <http://www.gnu.org/licenses/>.
*/

module match_ram #(parameter wordsize = 16, parameter lines = 16) (
    input logic clk, reset, enable, read, write,
    input logic [lines-1:0] Match,
    inout logic [wordsize-1:0] RData
);

/***** Brief Description *******
 * First Created by Max Waugaman 2015
 *
 * match_ram contains the RAM used by the TLB. This RAM uses 
 * the match lines generated by the CAM as an address.
 ******************************/

// Create RAM
logic [wordsize-1:0] RAM[lines-1:0];
logic [$clog2(lines)-1:0] RAM_Adr;

// Create Address for RAM (update digital logic to use Match directly)
priority_encoder #(lines) pe(Match, RAM_Adr);

// Initialize RAM to 0
integer i;

// RAM Write
always_ff @(posedge clk)
  begin
    if(reset) begin
      for(i = 0; i < lines; i = i + 1) begin
        RAM[i] <= '0;
      end
    end else begin
      if (write & enable) begin
        // Word Write
        RAM[RAM_Adr] <= RData;
      end
    end
  end

// Create Read Output
assign RData = !write ? RAM[RAM_Adr] : 'bz;

endmodule // cam
