`ifndef _cfg_vh_
`define _cfg_vh_

//`define ECAHCES 1
`define PROFILE 1

`endif
